//======================================================================
//
// experimental_code.v
// -------------------
// Module for testing curve25519 sub functions.
//
//
// Author: Joachim Strömbergson
// (c) 2015 Assured AB
//
//======================================================================


module experimental_code ();

  always @ init
    begin

    end

endmodule // experimental_code

//======================================================================
// EOF experimental_code.v
//======================================================================
